    Mac OS X            	   2  Y     �    TEXT                              ATTR      �   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     8   S  com.dropbox.attributes   [c\    e͋7     D?a*I9�XO��$�                                                      x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK��,��줪K�ܪ*G�������r[[���Z ՑP