    Mac OS X            	   2  Y     �    TEXT                              ATTR      �   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     8   S  com.dropbox.attributes   ��__    �"     D?a*I9�XO��$�                                                      x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%C�(WϜ4��bos�$o#�@_�t[[���Z ���