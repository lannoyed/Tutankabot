    Mac OS X            	   2   �                                           ATTR         �   X                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl   q��]    Tg�"     D?a*I9�XO��$�                                                      