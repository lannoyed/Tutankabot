    Mac OS X            	   2  Y     �                                      ATTR      �   �   �                  �     com.apple.lastuseddate#PS       �   H  com.apple.macl     8   S  com.dropbox.attributes   ���]    q	4     {�)��3NT��y�Tl� �1�EC����
�Ӧ�                                    x��VJ)�/Hʯ�O��I�L���ON�Q�R�V�ML����%����RK�%��H���r/W��D�,'w��0�|G[[���Z ��O